LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ctrl IS
  PORT